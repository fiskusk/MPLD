----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
----------------------------------------------------------------------------------
ENTITY TOP IS
  PORT(
    clk             : IN  STD_LOGIC;
    btn_i           : IN  STD_LOGIC_VECTOR (1 TO 4);
    sw_i            : IN  STD_LOGIC_VECTOR (1 TO 4);
    led_o           : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    disp_seg_o      : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    disp_dig_o      : OUT STD_LOGIC_VECTOR (4 DOWNTO 0)
  );
END TOP;
----------------------------------------------------------------------------------
ARCHITECTURE Structural OF TOP IS
----------------------------------------------------------------------------------


----------------------------------------------------------------------------------
BEGIN
----------------------------------------------------------------------------------


----------------------------------------------------------------------------------
END Structural;
----------------------------------------------------------------------------------
